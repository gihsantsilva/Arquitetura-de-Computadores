<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>1.76875,-2.6625,101.781,-54.2438</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>16,-8</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>19,-8</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>22,-8</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>25,-8</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>55,-8</position>
<input>
<ID>N_in2</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>59,-8</position>
<input>
<ID>N_in2</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>63,-8</position>
<input>
<ID>N_in2</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AI_XOR2</type>
<position>29.5,-14</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>29.5,-20.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>51,-28</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>51,-34</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>55,-6</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>59,-6</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>63,-6</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AE_OR2</type>
<position>60,-30.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>16,-6</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>19,-6</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>22,-6</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>25,-6</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AI_XOR3</type>
<position>41.5,-25</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_2</ID>17 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-21.5,25,-10</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-21.5 6</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-13,26.5,-13</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>25,-21.5,26.5,-21.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-15,19,-10</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-15,26.5,-15</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection>
<intersection>26.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>26.5,-19.5,26.5,-15</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-15 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-14,55,-9</points>
<connection>
<GID>10</GID>
<name>N_in2</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-14,55,-14</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-35,16,-10</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-35 1</intersection>
<intersection>-25 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-35,48,-35</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>16,-25,38.5,-25</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-29.5,57,-28</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54,-28,57,-28</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-34,57,-31.5</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54,-34,57,-34</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-30.5,63,-9</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32.5,-20.5,48,-20.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>36 4</intersection>
<intersection>48 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48,-29,48,-20.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>36,-23,36,-20.5</points>
<intersection>-23 5</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>36,-23,38.5,-23</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>36 4</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-33,22,-10</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-33 5</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-28.5,32,-28.5</points>
<intersection>22 0</intersection>
<intersection>32 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32,-28.5,32,-27</points>
<intersection>-28.5 1</intersection>
<intersection>-27 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>32,-27,38.5,-27</points>
<connection>
<GID>44</GID>
<name>IN_2</name></connection>
<intersection>32 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>22,-33,48,-33</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-25,59,-9</points>
<connection>
<GID>12</GID>
<name>N_in2</name></connection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-25,59,-25</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>48 2</intersection>
<intersection>59 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-27,48,-25</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-25 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 9></circuit>