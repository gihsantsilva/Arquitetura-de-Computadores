<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>1.39652,-4.06559,79.6441,-45.7153</PageViewport>
<gate>
<ID>4</ID>
<type>AA_AND3</type>
<position>52,-24</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>1 </input>
<input>
<ID>IN_2</ID>5 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_SMALL_INVERTER</type>
<position>39.5,-24</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>60,-24</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>20,-20</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>20,-24</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>20,-28</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41.5,-24,49,-24</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-24,59,-24</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-22,35.5,-20</points>
<intersection>-22 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-22,49,-22</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-20,35.5,-20</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-24,37.5,-24</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>6</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-28,49,-28</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>49 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49,-28,49,-26</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<intersection>-28 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 1>
<page 2>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 2>
<page 3>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 3>
<page 4>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 4>
<page 5>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 5>
<page 6>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 6>
<page 7>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 7>
<page 8>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 8>
<page 9>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 9></circuit>