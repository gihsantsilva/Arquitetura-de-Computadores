<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>1.74817,2.19848,93.6518,-43.2278</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>8,-5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>12,-5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>16,-5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>20,-5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>64,-5</position>
<input>
<ID>N_in2</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>68,-5</position>
<input>
<ID>N_in2</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>72,-5</position>
<input>
<ID>N_in2</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>76,-5</position>
<input>
<ID>N_in2</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>8,-2.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>12,-2.5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>16,-2.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>20,-2.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_AND2</type>
<position>27,-10</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_AND2</type>
<position>27,-16</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND2</type>
<position>27,-22</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_AND2</type>
<position>27,-28</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>AI_XOR2</type>
<position>43,-14.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_AND2</type>
<position>41.5,-23</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AI_XOR2</type>
<position>59.5,-24</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>64,-2.5</position>
<gparam>LABEL_TEXT R4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>69,-6.5</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>76,-2.5</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>72,-2.5</position>
<gparam>LABEL_TEXT R2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>73,-6.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>65,-6.5</position>
<gparam>LABEL_TEXT 8</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>77.5,-6.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>68,-2.5</position>
<gparam>LABEL_TEXT R3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_AND2</type>
<position>51.5,-31</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-11,8,-7</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-11,24,-11</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>8 0</intersection>
<intersection>24 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>24,-15,24,-11</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-11 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-9,16,-7</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-9,24,-9</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection>
<intersection>24 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>24,-23,24,-9</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>-9 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-17,20,-7</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-17,24,-17</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>20 0</intersection>
<intersection>24 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>24,-29,24,-17</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>-17 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-21,12,-7</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-21,24,-21</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>12 0</intersection>
<intersection>24 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>24,-27,24,-21</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-10,76,-6</points>
<connection>
<GID>16</GID>
<name>N_in2</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-10,76,-10</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-24,37,-13.5</points>
<intersection>-24 6</intersection>
<intersection>-22 5</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-13.5,40,-13.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>30 7</intersection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>37,-22,38.5,-22</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>37,-24,38.5,-24</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>30,-16,30,-13.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>-13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-22,37,-15.5</points>
<intersection>-22 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-15.5,40,-15.5</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-22,37,-22</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-14.5,72,-6</points>
<connection>
<GID>14</GID>
<name>N_in2</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-14.5,72,-14.5</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-23,56.5,-23</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>48.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>48.5,-30,48.5,-23</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-23 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-28,56.5,-28</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>48.5 7</intersection>
<intersection>56.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>56.5,-28,56.5,-25</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>48.5,-32,48.5,-28</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>-28 1</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-24,68,-6</points>
<connection>
<GID>12</GID>
<name>N_in2</name></connection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-24,68,-24</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-31,64,-6</points>
<connection>
<GID>10</GID>
<name>N_in2</name></connection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-31,64,-31</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>